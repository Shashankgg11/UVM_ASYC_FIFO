class afifo_wdriver extends uvm_driver #(afifo_seq_item);

	virtual afifo_if wvif;
	afifo_seq_item seq;

    `uvm_component_utils(afifo_wdriver)

    function new(string name = "afifo_wdriver", uvm_component parent);
		super.new(name, parent);
	endfunction

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
        if(!uvm_config_db #(virtual afifo_if)::get(this,"","vif",wvif))`uvm_error(get_type_name(), $sformatf("Failed to get WVIF"))
	endfunction

	virtual task run_phase(uvm_phase phase);
		forever 
		begin
			seq_item_port.get_next_item(seq);
			drive();
			seq_item_port.item_done();
		end
	endtask

	virtual task drive();
      repeat(1) @(wvif.wdriver_cb);
		wvif.wdata <= seq.wdata;
		wvif.winc <= seq.winc;
      `uvm_info(get_type_name(), $sformatf("Write_Driver DRIVER sent to DUT:, wdata = %0d, winc = %0d", wvif.wdata, wvif.winc), UVM_MEDIUM)
	endtask
endclass
